module InsFetch(oins, oadder, ohit, );



endmodule // main
